import lc3b_types::*

module test_tb

timeunit 1;
timeprecision ns;


blender dut
(

);


endmodule
