//####################################################################
//####################################################################
//####################################################################
//################ Created by Nick Moore  ############################
//################  for MP2 in ECE 411 at ############################
//################ University of Illinois ############################
//################ Fall 2015              ############################
//####################################################################
//####################################################################
//####################################################################
//#                                                                  #
//#   cache_datapath.sv                                              #
//#     Implements the datapath module for the LC3B cache            #
//#     controlled by the control module for the LC3B cache          #
//#     instantiate both in cache.sv and connect the inputs/outputs  #
//#                                                                  #
//####################################################################

import lc3b_types::*;

module cache_datapath
(
	//signals between cache and cpu datapath
	input lc3b_word mem_address,
	input lc3b_word mem_wdata,
	input [1:0] mem_byte_enable,
	output lc3b_word mem_rdata,

	//signals between cache and physical memory
	input cache_line pmem_rdata,
	output cache_line pmem_wdata,

	//signals between cache datapath and cache controller
	input clk,
	input valid_data,
	input dirty_data,
	input write1, write0,
	input pmem_wdatamux_sel,		//mux selects
	input datainmux1_sel, datainmux0_sel,	//mux selects
	output logic isValid1, isValid0,
	output logic isHit1, isHit0,		//logic determining if there was a hit
	output logic isDirty1, isDirty0,
	output cache_index index_out,
	output cache_tag tag_out,
	output cache_tag [1:0] tags,
	output cache_offset offset_out
);

//#############################################################################################################
//#############################################################################################################
//#############################################################################################################
//############################                                                 ################################
//############################                                                 ################################
//############################                 Variable Declarations           ################################
//############################                                                 ################################
//############################                                                 ################################
//############################                                                 ################################
//#############################################################################################################
//#############################################################################################################
//#############################################################################################################

cache_index index;				//set select stripped off of mem_address
cache_offset offset;				//word select stripped off of mem_address
cache_tag tag;					//set tag stripped off of mem_address
cache_line datainmux1_out, datainmux0_out;	//logic entering set ways
cache_line way1_out, way0_out;			//logic exiting set ways
cache_tag tag1_out, tag0_out;			//logic outputs from tag arrays
cache_line dataoutmux_out;			//connects dataoutmux to wordselectmux
cache_line blender1_out, blender0_out;		//outputs from the blenders to the datainmuxes


logic valid1_out, valid0_out;		//logic outputs from valid arrays
logic tagcompare1_out, tagcompare0_out;	//logic checking for tag hits
logic hitcheck1, hitcheck0;		//logic determining if each array has a hit
logic [7:0] decoder1_out, decoder0_out;	//logic from decoder as mux select lines in blender

logic dataoutmux_sel;			//select line from dataoutmux -- controlled by combinational logic

//#############################################################################################################
//#############################################################################################################
//#############################################################################################################
//############################                                                 ################################
//############################                                                 ################################
//############################               Variable Definitions              ################################
//############################                                                 ################################
//############################                                                 ################################
//############################                                                 ################################
//#############################################################################################################
//#############################################################################################################
//#############################################################################################################

assign isValid1 = valid1_out;
assign isValid0 = valid0_out;
assign index = mem_address[6:4];
assign index_out = index;
assign offset = mem_address[3:1];
assign tag = mem_address[15:7];
assign tag_out = tag;
assign isHit1 = hitcheck1;
assign isHit0 = hitcheck0;
assign hitcheck1 = valid1_out & tagcompare1_out;
assign hitcheck0 = valid0_out & tagcompare0_out;
assign dataoutmux_sel = hitcheck1;
assign tags[1] = tag1_out;
assign tags[0] = tag0_out;
assign offset_out = offset;

//#############################################################################################################
//#############################################################################################################
//#############################################################################################################
//############################                                                 ################################
//############################                                                 ################################
//############################              Associativity Ways                 ################################
//############################                                                 ################################
//############################                                                 ################################
//############################                                                 ################################
//#############################################################################################################
//#############################################################################################################
//#############################################################################################################

array way1 
(
    .clk(clk),
    .write(write1),
    .index(index),
    .datain(datainmux1_out),
    .dataout(way1_out)
);

array way0
(
    .clk(clk),
    .write(write0),
    .index(index),
    .datain(datainmux0_out),
    .dataout(way0_out)
);

//#############################################################################################################
//#############################################################################################################
//#############################################################################################################
//############################                                                 ################################
//############################                                                 ################################
//############################               Tag Arrays                        ################################
//############################                                                 ################################
//############################                                                 ################################
//############################                                                 ################################
//#############################################################################################################
//#############################################################################################################
//#############################################################################################################

array #(.width(9)) tag1
(
    .clk(clk),
    .write(write1),
    .index(index),
    .datain(tag),
    .dataout(tag1_out)
);

array #(.width(9)) tag0
(
    .clk(clk),
    .write(write0),
    .index(index),
    .datain(tag),
    .dataout(tag0_out)
);

compare tagcompare0
(
	.tag_a(tag0_out),
	.tag_b(tag),
	.isEqual(tagcompare0_out)
);

compare tagcompare1
(
	.tag_a(tag1_out),
	.tag_b(tag),
	.isEqual(tagcompare1_out)
);

//#############################################################################################################
//#############################################################################################################
//#############################################################################################################
//############################                                                 ################################
//############################                                                 ################################
//############################               Validity Check Arrays             ################################
//############################                                                 ################################
//############################                                                 ################################
//############################                                                 ################################
//#############################################################################################################
//#############################################################################################################
//#############################################################################################################

array #(.width(1)) valid1
(
    .clk(clk),
    .write(write1),
    .index(index),
    .datain(valid_data),
    .dataout(valid1_out)
);

array #(.width(1)) valid0
(
    .clk(clk),
    .write(write0),
    .index(index),
    .datain(valid_data),
    .dataout(valid0_out)
);

//#############################################################################################################
//#############################################################################################################
//#############################################################################################################
//############################                                                 ################################
//############################                                                 ################################
//############################               Dirty Bit Arrays                  ################################
//############################                                                 ################################
//############################                                                 ################################
//############################                                                 ################################
//#############################################################################################################
//#############################################################################################################
//#############################################################################################################

array #(.width(1)) dirty1
(
    .clk(clk),
    .write(write1),
    .index(index),
    .datain(dirty_data),
    .dataout(isDirty1)
);

array #(.width(1)) dirty0
(
    .clk(clk),
    .write(write0),
    .index(index),
    .datain(dirty_data),
    .dataout(isDirty0)
);

//#############################################################################################################
//#############################################################################################################
//#############################################################################################################
//############################                                                 ################################
//############################                                                 ################################
//############################                  Multiplexors                   ################################
//############################                                                 ################################
//############################                                                 ################################
//############################                                                 ################################
//#############################################################################################################
//#############################################################################################################
//#############################################################################################################

mux2 #(.width(128)) dataoutmux
(
	.a(way0_out),
	.b(way1_out),
	.sel(dataoutmux_sel),
	.f(dataoutmux_out)
);

mux8  wordselectmux
(
	.a(dataoutmux_out[0]),
	.b(dataoutmux_out[1]),
	.c(dataoutmux_out[2]),
	.d(dataoutmux_out[3]),
	.e(dataoutmux_out[4]),
	.f(dataoutmux_out[5]),
	.g(dataoutmux_out[6]),
	.h(dataoutmux_out[7]),
	.sel(offset),
	.i(mem_rdata)
);

mux2 #(.width(128)) pmem_wdatamux
(
	.a(way0_out),
	.b(way1_out),
	.sel(pmem_wdatamux_sel),
	.f(pmem_wdata)
);

mux2 #(.width(128)) datainmux1
(
	.a(blender1_out),
	.b(pmem_rdata),
	.sel(datainmux1_sel),
	.f(datainmux1_out)
);

mux2 #(.width(128)) datainmux0
(
	.a(blender0_out),
	.b(pmem_rdata),
	.sel(datainmux0_sel),
	.f(datainmux0_out)
);

//#############################################################################################################
//#############################################################################################################
//#############################################################################################################
//############################                                                 ################################
//############################                                                 ################################
//############################                     Blender                     ################################
//############################                (made from multiplexors)         ################################
//############################                                                 ################################
//############################                                                 ################################
//#############################################################################################################
//#############################################################################################################
//#############################################################################################################

blender blender0
(
	.in_line(way0_out),
	.offset(offset),
	.mem_byte_enable(mem_byte_enable),
	.data(mem_wdata),
	.out_line(blender0_out)
);

blender blender1
(
	.in_line(way1_out),
	.offset(offset),
	.mem_byte_enable(mem_byte_enable),
	.data(mem_wdata),
	.out_line(blender1_out)
);

endmodule : cache_datapath
