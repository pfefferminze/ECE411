module adder #(parameter width = 16)
(
	input logic [width - 1:0] a,b,
	output logic [width - 1:0] sum
);
assign sum = a + b;

endmodule : adder
