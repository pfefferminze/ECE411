import lc3b_types::*;
import cache_types::*;

module lru_tb;


   timeunit 1ns;
   timeprecision 1ps;

   logic [7:0] hit;
   logic 	   mem_resp;
   logic [1:0] out;
   logic 	   clk;
   logic [3:0][1:0] internals;
   

   initial clk = 0;
   always #1 clk = !clk;
   
   victim_lru dut(.*,.out(out));

   initial begin : waveform_generation
	  hit = 8'h1;
	  index = 3'h0;
	  mem_resp = 0;
	  $display("initial out = %d",out);
	  #5 mem_resp = 1;
	  $display("initial out = %d",out);
	  #5 mem_resp = 0;
	  hit = 8'h2;
	  $display("initial out = %d",out);
	  #5 mem_resp = 1;
	  $display("initial out = %d",out);
	  #5 mem_resp = 0;
	  hit = 8'h4;
	  $display("initial out = %d",out);
	  #5 mem_resp = 1;
	  $display("initial out = %d",out);
	  #5 mem_resp = 0;
	  hit = 8'h8;
	  $display("initial out = %d",out);
	  #5 mem_resp = 1;
	  $display("initial out = %d",out);
	  #5 mem_resp = 0;
	  hit = 8'h10;
	  $display("initial out = %d",out);
	  #5 mem_resp = 1;
	  $display("initial out = %d",out);
	  #5 mem_resp = 0;
	  hit = 8'h20;
	  $display("initial out = %d",out);
	  #5 mem_resp = 1;
	  $display("initial out = %d",out);
	  #5 mem_resp = 0;
	  hit = 8'h40;
	  $display("initial out = %d",out);
	  #5 mem_resp = 1;
	  $display("initial out = %d",out);
	  #5 mem_resp = 0;
	  hit = 8'h80;
	  $display("initial out = %d",out);
	  #5 mem_resp = 1;
	  $display("initial out = %d",out);
	  #5 mem_resp = 0;
	  hit = 8'h0;
	  $display("initial out = %d",out);
	  #5 mem_resp = 1;
	  $display("initial out = %d",out);
	  #5 mem_resp = 0;
	  hit = 8'h4;
	  $display("initial out = %d",out);
	  #5 mem_resp = 1;
	  $display("initial out = %d",out);
	  #5 mem_resp = 0;
	  hit = 8'h2;
	  $display("initial out = %d",out);
	  #5 mem_resp = 1;
	  $display("initial out = %d",out);
	  #5 mem_resp = 0;
	  hit = 8'h2;
	  $display("initial out = %d",out);
	  #5 mem_resp = 1;
	  $display("initial out = %d",out);
	  #5 mem_resp = 0;
	  hit = 8'h1;
	  $display("out = %d",out);
	  #5 mem_resp=1;
	  $display("out = %d",out);
	  #5
	  hit = 8'h1;
	  index = 3'h1;
	  mem_resp = 0;
	  $display("initial out = %d",out);
	  #5 mem_resp = 1;
	  $display("initial out = %d",out);
	  #5 mem_resp = 0;
	  hit = 8'h2;
	  $display("initial out = %d",out);
	  #5 mem_resp = 1;
	  $display("initial out = %d",out);
	  #5 mem_resp = 0;
	  hit = 8'h4;
	  $display("initial out = %d",out);
	  #5 mem_resp = 1;
	  $display("initial out = %d",out);
	  #5 mem_resp = 0;
	  hit = 8'h8;
	  $display("initial out = %d",out);
	  #5 mem_resp = 1;
	  $display("initial out = %d",out);
	  #5 mem_resp = 0;
	  hit = 8'h10;
	  $display("initial out = %d",out);
	  #5 mem_resp = 1;
	  $display("initial out = %d",out);
	  #5 mem_resp = 0;
	  hit = 8'h20;
	  $display("initial out = %d",out);
	  #5 mem_resp = 1;
	  $display("initial out = %d",out);
	  #5 mem_resp = 0;
	  hit = 8'h40;
	  $display("initial out = %d",out);
	  #5 mem_resp = 1;
	  $display("initial out = %d",out);
	  #5 mem_resp = 0;
	  hit = 8'h80;
	  $display("initial out = %d",out);
	  #5 mem_resp = 1;
	  $display("initial out = %d",out);
	  #5 mem_resp = 0;
	  hit = 8'h0;
	  $display("initial out = %d",out);
	  #5 mem_resp = 1;
	  $display("initial out = %d",out);
	  #5 mem_resp = 0;
	  hit = 8'h4;
	  $display("initial out = %d",out);
	  #5 mem_resp = 1;
	  $display("initial out = %d",out);
	  #5 mem_resp = 0;
	  hit = 8'h2;
	  $display("initial out = %d",out);
	  #5 mem_resp = 1;
	  $display("initial out = %d",out);
	  #5 mem_resp = 0;
	  hit = 8'h2;
	  $display("initial out = %d",out);
	  #5 mem_resp = 1;
	  $display("initial out = %d",out);
	  #5 mem_resp = 0;
	  hit = 8'h1;
	  $display("out = %d",out);
	  #5 mem_resp=1;
	  $display("out = %d",out);
	  #5
	  hit = 8'h1;
	  index = 3'h2;
	  mem_resp = 0;
	  $display("initial out = %d",out);
	  #5 mem_resp = 1;
	  $display("initial out = %d",out);
	  #5 mem_resp = 0;
	  hit = 8'h2;
	  $display("initial out = %d",out);
	  #5 mem_resp = 1;
	  $display("initial out = %d",out);
	  #5 mem_resp = 0;
	  hit = 8'h4;
	  $display("initial out = %d",out);
	  #5 mem_resp = 1;
	  $display("initial out = %d",out);
	  #5 mem_resp = 0;
	  hit = 8'h8;
	  $display("initial out = %d",out);
	  #5 mem_resp = 1;
	  $display("initial out = %d",out);
	  #5 mem_resp = 0;
	  hit = 8'h10;
	  $display("initial out = %d",out);
	  #5 mem_resp = 1;
	  $display("initial out = %d",out);
	  #5 mem_resp = 0;
	  hit = 8'h20;
	  $display("initial out = %d",out);
	  #5 mem_resp = 1;
	  $display("initial out = %d",out);
	  #5 mem_resp = 0;
	  hit = 8'h40;
	  $display("initial out = %d",out);
	  #5 mem_resp = 1;
	  $display("initial out = %d",out);
	  #5 mem_resp = 0;
	  hit = 8'h80;
	  $display("initial out = %d",out);
	  #5 mem_resp = 1;
	  $display("initial out = %d",out);
	  #5 mem_resp = 0;
	  hit = 8'h0;
	  $display("initial out = %d",out);
	  #5 mem_resp = 1;
	  $display("initial out = %d",out);
	  #5 mem_resp = 0;
	  hit = 8'h4;
	  $display("initial out = %d",out);
	  #5 mem_resp = 1;
	  $display("initial out = %d",out);
	  #5 mem_resp = 0;
	  hit = 8'h2;
	  $display("initial out = %d",out);
	  #5 mem_resp = 1;
	  $display("initial out = %d",out);
	  #5 mem_resp = 0;
	  hit = 8'h2;
	  $display("initial out = %d",out);
	  #5 mem_resp = 1;
	  $display("initial out = %d",out);
	  #5 mem_resp = 0;
	  hit = 8'h1;
	  $display("out = %d",out);
	  #5 mem_resp=1;
	  $display("out = %d",out);
	  
	  #5
	  hit = 8'h1;
	  index = 3'h3;
	  mem_resp = 0;
	  $display("initial out = %d",out);
	  #5 mem_resp = 1;
	  $display("initial out = %d",out);
	  #5 mem_resp = 0;
	  hit = 8'h2;
	  $display("initial out = %d",out);
	  #5 mem_resp = 1;
	  $display("initial out = %d",out);
	  #5 mem_resp = 0;
	  hit = 8'h4;
	  $display("initial out = %d",out);
	  #5 mem_resp = 1;
	  $display("initial out = %d",out);
	  #5 mem_resp = 0;
	  hit = 8'h8;
	  $display("initial out = %d",out);
	  #5 mem_resp = 1;
	  $display("initial out = %d",out);
	  #5 mem_resp = 0;
	  hit = 8'h10;
	  $display("initial out = %d",out);
	  #5 mem_resp = 1;
	  $display("initial out = %d",out);
	  #5 mem_resp = 0;
	  hit = 8'h20;
	  $display("initial out = %d",out);
	  #5 mem_resp = 1;
	  $display("initial out = %d",out);
	  #5 mem_resp = 0;
	  hit = 8'h40;
	  $display("initial out = %d",out);
	  #5 mem_resp = 1;
	  $display("initial out = %d",out);
	  #5 mem_resp = 0;
	  hit = 8'h80;
	  $display("initial out = %d",out);
	  #5 mem_resp = 1;
	  $display("initial out = %d",out);
	  #5 mem_resp = 0;
	  hit = 8'h0;
	  $display("initial out = %d",out);
	  #5 mem_resp = 1;
	  $display("initial out = %d",out);
	  #5 mem_resp = 0;
	  hit = 8'h4;
	  $display("initial out = %d",out);
	  #5 mem_resp = 1;
	  $display("initial out = %d",out);
	  #5 mem_resp = 0;
	  hit = 8'h2;
	  $display("initial out = %d",out);
	  #5 mem_resp = 1;
	  $display("initial out = %d",out);
	  #5 mem_resp = 0;
	  hit = 8'h2;
	  $display("initial out = %d",out);
	  #5 mem_resp = 1;
	  $display("initial out = %d",out);
	  #5 mem_resp = 0;
	  hit = 8'h1;
	  $display("out = %d",out);
	  #5 mem_resp=1;
	  $display("out = %d",out);

	  #5
	  hit = 8'h1;
	  index = 3'h4;
	  mem_resp = 0;
	  $display("initial out = %d",out);
	  #5 mem_resp = 1;
	  $display("initial out = %d",out);
	  #5 mem_resp = 0;
	  hit = 8'h2;
	  $display("initial out = %d",out);
	  #5 mem_resp = 1;
	  $display("initial out = %d",out);
	  #5 mem_resp = 0;
	  hit = 8'h4;
	  $display("initial out = %d",out);
	  #5 mem_resp = 1;
	  $display("initial out = %d",out);
	  #5 mem_resp = 0;
	  hit = 8'h8;
	  $display("initial out = %d",out);
	  #5 mem_resp = 1;
	  $display("initial out = %d",out);
	  #5 mem_resp = 0;
	  hit = 8'h10;
	  $display("initial out = %d",out);
	  #5 mem_resp = 1;
	  $display("initial out = %d",out);
	  #5 mem_resp = 0;
	  hit = 8'h20;
	  $display("initial out = %d",out);
	  #5 mem_resp = 1;
	  $display("initial out = %d",out);
	  #5 mem_resp = 0;
	  hit = 8'h40;
	  $display("initial out = %d",out);
	  #5 mem_resp = 1;
	  $display("initial out = %d",out);
	  #5 mem_resp = 0;
	  hit = 8'h80;
	  $display("initial out = %d",out);
	  #5 mem_resp = 1;
	  $display("initial out = %d",out);
	  #5 mem_resp = 0;
	  hit = 8'h0;
	  $display("initial out = %d",out);
	  #5 mem_resp = 1;
	  $display("initial out = %d",out);
	  #5 mem_resp = 0;
	  hit = 8'h4;
	  $display("initial out = %d",out);
	  #5 mem_resp = 1;
	  $display("initial out = %d",out);
	  #5 mem_resp = 0;
	  hit = 8'h2;
	  $display("initial out = %d",out);
	  #5 mem_resp = 1;
	  $display("initial out = %d",out);
	  #5 mem_resp = 0;
	  hit = 8'h2;
	  $display("initial out = %d",out);
	  #5 mem_resp = 1;
	  $display("initial out = %d",out);
	  #5 mem_resp = 0;
	  hit = 8'h1;
	  $display("out = %d",out);
	  #5 mem_resp=1;
	  $display("out = %d",out);

	  #5
	  hit = 8'h1;
	  index = 3'h5;
	  mem_resp = 0;
	  $display("initial out = %d",out);
	  #5 mem_resp = 1;
	  $display("initial out = %d",out);
	  #5 mem_resp = 0;
	  hit = 8'h2;
	  $display("initial out = %d",out);
	  #5 mem_resp = 1;
	  $display("initial out = %d",out);
	  #5 mem_resp = 0;
	  hit = 8'h4;
	  $display("initial out = %d",out);
	  #5 mem_resp = 1;
	  $display("initial out = %d",out);
	  #5 mem_resp = 0;
	  hit = 8'h8;
	  $display("initial out = %d",out);
	  #5 mem_resp = 1;
	  $display("initial out = %d",out);
	  #5 mem_resp = 0;
	  hit = 8'h10;
	  $display("initial out = %d",out);
	  #5 mem_resp = 1;
	  $display("initial out = %d",out);
	  #5 mem_resp = 0;
	  hit = 8'h20;
	  $display("initial out = %d",out);
	  #5 mem_resp = 1;
	  $display("initial out = %d",out);
	  #5 mem_resp = 0;
	  hit = 8'h40;
	  $display("initial out = %d",out);
	  #5 mem_resp = 1;
	  $display("initial out = %d",out);
	  #5 mem_resp = 0;
	  hit = 8'h80;
	  $display("initial out = %d",out);
	  #5 mem_resp = 1;
	  $display("initial out = %d",out);
	  #5 mem_resp = 0;
	  hit = 8'h0;
	  $display("initial out = %d",out);
	  #5 mem_resp = 1;
	  $display("initial out = %d",out);
	  #5 mem_resp = 0;
	  hit = 8'h4;
	  $display("initial out = %d",out);
	  #5 mem_resp = 1;
	  $display("initial out = %d",out);
	  #5 mem_resp = 0;
	  hit = 8'h2;
	  $display("initial out = %d",out);
	  #5 mem_resp = 1;
	  $display("initial out = %d",out);
	  #5 mem_resp = 0;
	  hit = 8'h2;
	  $display("initial out = %d",out);
	  #5 mem_resp = 1;
	  $display("initial out = %d",out);
	  #5 mem_resp = 0;
	  hit = 8'h1;
	  $display("out = %d",out);
	  #5 mem_resp=1;
	  $display("out = %d",out);

	  #5
	  hit = 8'h1;
	  index = 3'h6;
	  mem_resp = 0;
	  $display("initial out = %d",out);
	  #5 mem_resp = 1;
	  $display("initial out = %d",out);
	  #5 mem_resp = 0;
	  hit = 8'h2;
	  $display("initial out = %d",out);
	  #5 mem_resp = 1;
	  $display("initial out = %d",out);
	  #5 mem_resp = 0;
	  hit = 8'h4;
	  $display("initial out = %d",out);
	  #5 mem_resp = 1;
	  $display("initial out = %d",out);
	  #5 mem_resp = 0;
	  hit = 8'h8;
	  $display("initial out = %d",out);
	  #5 mem_resp = 1;
	  $display("initial out = %d",out);
	  #5 mem_resp = 0;
	  hit = 8'h10;
	  $display("initial out = %d",out);
	  #5 mem_resp = 1;
	  $display("initial out = %d",out);
	  #5 mem_resp = 0;
	  hit = 8'h20;
	  $display("initial out = %d",out);
	  #5 mem_resp = 1;
	  $display("initial out = %d",out);
	  #5 mem_resp = 0;
	  hit = 8'h40;
	  $display("initial out = %d",out);
	  #5 mem_resp = 1;
	  $display("initial out = %d",out);
	  #5 mem_resp = 0;
	  hit = 8'h80;
	  $display("initial out = %d",out);
	  #5 mem_resp = 1;
	  $display("initial out = %d",out);
	  #5 mem_resp = 0;
	  hit = 8'h0;
	  $display("initial out = %d",out);
	  #5 mem_resp = 1;
	  $display("initial out = %d",out);
	  #5 mem_resp = 0;
	  hit = 8'h4;
	  $display("initial out = %d",out);
	  #5 mem_resp = 1;
	  $display("initial out = %d",out);
	  #5 mem_resp = 0;
	  hit = 8'h2;
	  $display("initial out = %d",out);
	  #5 mem_resp = 1;
	  $display("initial out = %d",out);
	  #5 mem_resp = 0;
	  hit = 8'h2;
	  $display("initial out = %d",out);
	  #5 mem_resp = 1;
	  $display("initial out = %d",out);
	  #5 mem_resp = 0;
	  hit = 8'h1;
	  $display("out = %d",out);
	  #5 mem_resp=1;
	  $display("out = %d",out);

	  #5
	  hit = 8'h1;
	  index = 3'h7;
	  mem_resp = 0;
	  $display("initial out = %d",out);
	  #5 mem_resp = 1;
	  $display("initial out = %d",out);
	  #5 mem_resp = 0;
	  hit = 8'h2;
	  $display("initial out = %d",out);
	  #5 mem_resp = 1;
	  $display("initial out = %d",out);
	  #5 mem_resp = 0;
	  hit = 8'h4;
	  $display("initial out = %d",out);
	  #5 mem_resp = 1;
	  $display("initial out = %d",out);
	  #5 mem_resp = 0;
	  hit = 8'h8;
	  $display("initial out = %d",out);
	  #5 mem_resp = 1;
	  $display("initial out = %d",out);
	  #5 mem_resp = 0;
	  hit = 8'h10;
	  $display("initial out = %d",out);
	  #5 mem_resp = 1;
	  $display("initial out = %d",out);
	  #5 mem_resp = 0;
	  hit = 8'h20;
	  $display("initial out = %d",out);
	  #5 mem_resp = 1;
	  $display("initial out = %d",out);
	  #5 mem_resp = 0;
	  hit = 8'h40;
	  $display("initial out = %d",out);
	  #5 mem_resp = 1;
	  $display("initial out = %d",out);
	  #5 mem_resp = 0;
	  hit = 8'h80;
	  $display("initial out = %d",out);
	  #5 mem_resp = 1;
	  $display("initial out = %d",out);
	  #5 mem_resp = 0;
	  hit = 8'h0;
	  $display("initial out = %d",out);
	  #5 mem_resp = 1;
	  $display("initial out = %d",out);
	  #5 mem_resp = 0;
	  hit = 8'h4;
	  $display("initial out = %d",out);
	  #5 mem_resp = 1;
	  $display("initial out = %d",out);
	  #5 mem_resp = 0;
	  hit = 8'h2;
	  $display("initial out = %d",out);
	  #5 mem_resp = 1;
	  $display("initial out = %d",out);
	  #5 mem_resp = 0;
	  hit = 8'h2;
	  $display("initial out = %d",out);
	  #5 mem_resp = 1;
	  $display("initial out = %d",out);
	  #5 mem_resp = 0;
	  hit = 8'h1;
	  $display("out = %d",out);
	  #5 mem_resp=1;
	  $display("out = %d",out);

	  #5
	  hit = 8'h1;
	  index = 3'h0;
	  mem_resp = 0;
	  $display("initial out = %d",out);
	  #5 mem_resp = 1;
	  $display("initial out = %d",out);
	  #5 mem_resp = 0;
	  hit = 8'h2;
	  $display("initial out = %d",out);
	  #5 mem_resp = 1;
	  $display("initial out = %d",out);
	  #5 mem_resp = 0;
	  hit = 8'h4;
	  $display("initial out = %d",out);
	  #5 mem_resp = 1;
	  $display("initial out = %d",out);
	  #5 mem_resp = 0;
	  hit = 8'h8;
	  $display("initial out = %d",out);
	  #5 mem_resp = 1;
	  $display("initial out = %d",out);
	  #5 mem_resp = 0;
	  hit = 8'h10;
	  $display("initial out = %d",out);
	  #5 mem_resp = 1;
	  $display("initial out = %d",out);
	  #5 mem_resp = 0;
	  hit = 8'h20;
	  $display("initial out = %d",out);
	  #5 mem_resp = 1;
	  $display("initial out = %d",out);
	  #5 mem_resp = 0;
	  hit = 8'h40;
	  $display("initial out = %d",out);
	  #5 mem_resp = 1;
	  $display("initial out = %d",out);
	  #5 mem_resp = 0;
	  hit = 8'h80;
	  $display("initial out = %d",out);
	  #5 mem_resp = 1;
	  $display("initial out = %d",out);
	  #5 mem_resp = 0;
	  hit = 8'h0;
	  $display("initial out = %d",out);
	  #5 mem_resp = 1;
	  $display("initial out = %d",out);
	  #5 mem_resp = 0;
	  hit = 8'h4;
	  $display("initial out = %d",out);
	  #5 mem_resp = 1;
	  $display("initial out = %d",out);
	  #5 mem_resp = 0;
	  hit = 8'h2;
	  $display("initial out = %d",out);
	  #5 mem_resp = 1;
	  $display("initial out = %d",out);
	  #5 mem_resp = 0;
	  hit = 8'h2;
	  $display("initial out = %d",out);
	  #5 mem_resp = 1;
	  $display("initial out = %d",out);
	  #5 mem_resp = 0;
	  hit = 8'h1;
	  $display("out = %d",out);
	  #5 mem_resp=1;
	  $display("out = %d",out);

	  #5
	  hit = 8'h1;
	  index = 3'h1;
	  mem_resp = 0;
	  $display("initial out = %d",out);
	  #5 mem_resp = 1;
	  $display("initial out = %d",out);
	  #5 mem_resp = 0;
	  hit = 8'h2;
	  $display("initial out = %d",out);
	  #5 mem_resp = 1;
	  $display("initial out = %d",out);
	  #5 mem_resp = 0;
	  hit = 8'h4;
	  $display("initial out = %d",out);
	  #5 mem_resp = 1;
	  $display("initial out = %d",out);
	  #5 mem_resp = 0;
	  hit = 8'h8;
	  $display("initial out = %d",out);
	  #5 mem_resp = 1;
	  $display("initial out = %d",out);
	  #5 mem_resp = 0;
	  hit = 8'h10;
	  $display("initial out = %d",out);
	  #5 mem_resp = 1;
	  $display("initial out = %d",out);
	  #5 mem_resp = 0;
	  hit = 8'h20;
	  $display("initial out = %d",out);
	  #5 mem_resp = 1;
	  $display("initial out = %d",out);
	  #5 mem_resp = 0;
	  hit = 8'h40;
	  $display("initial out = %d",out);
	  #5 mem_resp = 1;
	  $display("initial out = %d",out);
	  #5 mem_resp = 0;
	  hit = 8'h80;
	  $display("initial out = %d",out);
	  #5 mem_resp = 1;
	  $display("initial out = %d",out);
	  #5 mem_resp = 0;
	  hit = 8'h0;
	  $display("initial out = %d",out);
	  #5 mem_resp = 1;
	  $display("initial out = %d",out);
	  #5 mem_resp = 0;
	  hit = 8'h4;
	  $display("initial out = %d",out);
	  #5 mem_resp = 1;
	  $display("initial out = %d",out);
	  #5 mem_resp = 0;
	  hit = 8'h2;
	  $display("initial out = %d",out);
	  #5 mem_resp = 1;
	  $display("initial out = %d",out);
	  #5 mem_resp = 0;
	  hit = 8'h2;
	  $display("initial out = %d",out);
	  #5 mem_resp = 1;
	  $display("initial out = %d",out);
	  #5 mem_resp = 0;
	  hit = 8'h1;
	  $display("out = %d",out);
	  #5 mem_resp=1;
	  $display("out = %d",out);
   end : waveform_generation

endmodule // lru_tb
