import lc3b_types::*;
import cache_types::*;

module victim_lru_tb;


   timeunit 1ns;
   timeprecision 1ps;
   logic [1:0] out;
   logic [3:0] hit;
   logic 	   mem_resp;
   logic [1:0] l_r_u;
   logic 	   clk;
   logic [3:0][1:0] internals;
   

   initial clk = 0;
   always #1 clk = !clk;
   
   victim_lru dut(.*);

   initial begin : waveform_generation
	  hit = 4'h1;
	  mem_resp = 0;
	  $display("initial l_r_u = %d",l_r_u);
	  #5 mem_resp = 1;
	  $display("initial l_r_u = %d",l_r_u);
	  #5 mem_resp = 0;
	  hit = 4'h2;
	  $display("initial l_r_u = %d",l_r_u);
	  #5 mem_resp = 1;
	  $display("initial l_r_u = %d",l_r_u);
	  #5 mem_resp = 0;
	  hit = 4'h4;
	  $display("initial l_r_u = %d",l_r_u);
	  #5 mem_resp = 1;
	  $display("initial l_r_u = %d",l_r_u);
	  #5 mem_resp = 0;
	  hit = 4'h8;
	  $display("initial l_r_u = %d",l_r_u);
	  #5 mem_resp = 1;
	  $display("initial l_r_u = %d",l_r_u);
	  #5 mem_resp = 0;
	  hit = 4'h1;
	  $display("initial l_r_u = %d",l_r_u);
	  #5 mem_resp = 1;
	  $display("initial l_r_u = %d",l_r_u);
	  #5 mem_resp = 0;
	  hit = 4'h2;
	  $display("initial l_r_u = %d",l_r_u);
	  #5 mem_resp = 1;
	  $display("initial l_r_u = %d",l_r_u);
	  #5 mem_resp = 0;
	  hit = 4'h4;
	  $display("initial l_r_u = %d",l_r_u);
	  #5 mem_resp = 1;
	  $display("initial l_r_u = %d",l_r_u);
	  #5 mem_resp = 0;
	  hit = 4'h8;
	  $display("initial l_r_u = %d",l_r_u);
	  #5 mem_resp = 1;
	  $display("initial l_r_u = %d",l_r_u);
	  #5 mem_resp = 0;
	  hit = 4'h0;
	  $display("initial l_r_u = %d",l_r_u);
	  #5 mem_resp = 1;
	  $display("initial l_r_u = %d",l_r_u);
	  #5 mem_resp = 0;
	  hit = 4'h4;
	  $display("initial l_r_u = %d",l_r_u);
	  #5 mem_resp = 1;
	  $display("initial l_r_u = %d",l_r_u);
	  #5 mem_resp = 0;
	  hit = 4'h2;
	  $display("initial l_r_u = %d",l_r_u);
	  #5 mem_resp = 1;
	  $display("initial l_r_u = %d",l_r_u);
	  #5 mem_resp = 0;
	  hit = 4'h2;
	  $display("initial l_r_u = %d",l_r_u);
	  #5 mem_resp = 1;
	  $display("initial l_r_u = %d",l_r_u);
	  #5 mem_resp = 0;
	  hit = 4'h1;
	  $display("l_r_u = %d",l_r_u);
	  #5 mem_resp=1;
	  $display("l_r_u = %d",l_r_u);
	  #5
	  hit = 4'h1;
	  mem_resp = 0;
	  $display("initial l_r_u = %d",l_r_u);
	  #5 mem_resp = 1;
	  $display("initial l_r_u = %d",l_r_u);
	  #5 mem_resp = 0;
	  hit = 4'h2;
	  $display("initial l_r_u = %d",l_r_u);
	  #5 mem_resp = 1;
	  $display("initial l_r_u = %d",l_r_u);
	  #5 mem_resp = 0;
	  hit = 4'h4;
	  $display("initial l_r_u = %d",l_r_u);
	  #5 mem_resp = 1;
	  $display("initial l_r_u = %d",l_r_u);
	  #5 mem_resp = 0;
	  hit = 4'h8;
	  $display("initial l_r_u = %d",l_r_u);
	  #5 mem_resp = 1;
	  $display("initial l_r_u = %d",l_r_u);
	  #5 mem_resp = 0;
	  hit = 4'h1;
	  $display("initial l_r_u = %d",l_r_u);
	  #5 mem_resp = 1;
	  $display("initial l_r_u = %d",l_r_u);
	  #5 mem_resp = 0;
	  hit = 4'h2;
	  $display("initial l_r_u = %d",l_r_u);
	  #5 mem_resp = 1;
	  $display("initial l_r_u = %d",l_r_u);
	  #5 mem_resp = 0;
	  hit = 4'h4;
	  $display("initial l_r_u = %d",l_r_u);
	  #5 mem_resp = 1;
	  $display("initial l_r_u = %d",l_r_u);
	  #5 mem_resp = 0;
	  hit = 4'h8;
	  $display("initial l_r_u = %d",l_r_u);
	  #5 mem_resp = 1;
	  $display("initial l_r_u = %d",l_r_u);
	  #5 mem_resp = 0;
	  hit = 4'h0;
	  $display("initial l_r_u = %d",l_r_u);
	  #5 mem_resp = 1;
	  $display("initial l_r_u = %d",l_r_u);
	  #5 mem_resp = 0;
	  hit = 4'h4;
	  $display("initial l_r_u = %d",l_r_u);
	  #5 mem_resp = 1;
	  $display("initial l_r_u = %d",l_r_u);
	  #5 mem_resp = 0;
	  hit = 4'h2;
	  $display("initial l_r_u = %d",l_r_u);
	  #5 mem_resp = 1;
	  $display("initial l_r_u = %d",l_r_u);
	  #5 mem_resp = 0;
	  hit = 4'h2;
	  $display("initial l_r_u = %d",l_r_u);
	  #5 mem_resp = 1;
	  $display("initial l_r_u = %d",l_r_u);
	  #5 mem_resp = 0;
	  hit = 4'h1;
	  $display("l_r_u = %d",l_r_u);
	  #5 mem_resp=1;
	  $display("l_r_u = %d",l_r_u);
	  #5
	  hit = 4'h1;
	  mem_resp = 0;
	  $display("initial l_r_u = %d",l_r_u);
	  #5 mem_resp = 1;
	  $display("initial l_r_u = %d",l_r_u);
	  #5 mem_resp = 0;
	  hit = 4'h2;
	  $display("initial l_r_u = %d",l_r_u);
	  #5 mem_resp = 1;
	  $display("initial l_r_u = %d",l_r_u);
	  #5 mem_resp = 0;
	  hit = 4'h4;
	  $display("initial l_r_u = %d",l_r_u);
	  #5 mem_resp = 1;
	  $display("initial l_r_u = %d",l_r_u);
	  #5 mem_resp = 0;
	  hit = 4'h8;
	  $display("initial l_r_u = %d",l_r_u);
	  #5 mem_resp = 1;
	  $display("initial l_r_u = %d",l_r_u);
	  #5 mem_resp = 0;
	  hit = 4'h1;
	  $display("initial l_r_u = %d",l_r_u);
	  #5 mem_resp = 1;
	  $display("initial l_r_u = %d",l_r_u);
	  #5 mem_resp = 0;
	  hit = 4'h2;
	  $display("initial l_r_u = %d",l_r_u);
	  #5 mem_resp = 1;
	  $display("initial l_r_u = %d",l_r_u);
	  #5 mem_resp = 0;
	  hit = 4'h4;
	  $display("initial l_r_u = %d",l_r_u);
	  #5 mem_resp = 1;
	  $display("initial l_r_u = %d",l_r_u);
	  #5 mem_resp = 0;
	  hit = 4'h8;
	  $display("initial l_r_u = %d",l_r_u);
	  #5 mem_resp = 1;
	  $display("initial l_r_u = %d",l_r_u);
	  #5 mem_resp = 0;
	  hit = 4'h0;
	  $display("initial l_r_u = %d",l_r_u);
	  #5 mem_resp = 1;
	  $display("initial l_r_u = %d",l_r_u);
	  #5 mem_resp = 0;
	  hit = 4'h4;
	  $display("initial l_r_u = %d",l_r_u);
	  #5 mem_resp = 1;
	  $display("initial l_r_u = %d",l_r_u);
	  #5 mem_resp = 0;
	  hit = 4'h2;
	  $display("initial l_r_u = %d",l_r_u);
	  #5 mem_resp = 1;
	  $display("initial l_r_u = %d",l_r_u);
	  #5 mem_resp = 0;
	  hit = 4'h2;
	  $display("initial l_r_u = %d",l_r_u);
	  #5 mem_resp = 1;
	  $display("initial l_r_u = %d",l_r_u);
	  #5 mem_resp = 0;
	  hit = 4'h1;
	  $display("l_r_u = %d",l_r_u);
	  #5 mem_resp=1;
	  $display("l_r_u = %d",l_r_u);
	  
	  #5
	  hit = 4'h1;
	  mem_resp = 0;
	  $display("initial l_r_u = %d",l_r_u);
	  #5 mem_resp = 1;
	  $display("initial l_r_u = %d",l_r_u);
	  #5 mem_resp = 0;
	  hit = 4'h2;
	  $display("initial l_r_u = %d",l_r_u);
	  #5 mem_resp = 1;
	  $display("initial l_r_u = %d",l_r_u);
	  #5 mem_resp = 0;
	  hit = 4'h4;
	  $display("initial l_r_u = %d",l_r_u);
	  #5 mem_resp = 1;
	  $display("initial l_r_u = %d",l_r_u);
	  #5 mem_resp = 0;
	  hit = 4'h8;
	  $display("initial l_r_u = %d",l_r_u);
	  #5 mem_resp = 1;
	  $display("initial l_r_u = %d",l_r_u);
	  #5 mem_resp = 0;
	  hit = 4'h1;
	  $display("initial l_r_u = %d",l_r_u);
	  #5 mem_resp = 1;
	  $display("initial l_r_u = %d",l_r_u);
	  #5 mem_resp = 0;
	  hit = 4'h2;
	  $display("initial l_r_u = %d",l_r_u);
	  #5 mem_resp = 1;
	  $display("initial l_r_u = %d",l_r_u);
	  #5 mem_resp = 0;
	  hit = 4'h4;
	  $display("initial l_r_u = %d",l_r_u);
	  #5 mem_resp = 1;
	  $display("initial l_r_u = %d",l_r_u);
	  #5 mem_resp = 0;
	  hit = 4'h8;
	  $display("initial l_r_u = %d",l_r_u);
	  #5 mem_resp = 1;
	  $display("initial l_r_u = %d",l_r_u);
	  #5 mem_resp = 0;
	  hit = 4'h0;
	  $display("initial l_r_u = %d",l_r_u);
	  #5 mem_resp = 1;
	  $display("initial l_r_u = %d",l_r_u);
	  #5 mem_resp = 0;
	  hit = 4'h4;
	  $display("initial l_r_u = %d",l_r_u);
	  #5 mem_resp = 1;
	  $display("initial l_r_u = %d",l_r_u);
	  #5 mem_resp = 0;
	  hit = 4'h2;
	  $display("initial l_r_u = %d",l_r_u);
	  #5 mem_resp = 1;
	  $display("initial l_r_u = %d",l_r_u);
	  #5 mem_resp = 0;
	  hit = 4'h2;
	  $display("initial l_r_u = %d",l_r_u);
	  #5 mem_resp = 1;
	  $display("initial l_r_u = %d",l_r_u);
	  #5 mem_resp = 0;
	  hit = 4'h1;
	  $display("l_r_u = %d",l_r_u);
	  #5 mem_resp=1;
	  $display("l_r_u = %d",l_r_u);

	  #5
	  hit = 4'h1;
	  mem_resp = 0;
	  $display("initial l_r_u = %d",l_r_u);
	  #5 mem_resp = 1;
	  $display("initial l_r_u = %d",l_r_u);
	  #5 mem_resp = 0;
	  hit = 4'h2;
	  $display("initial l_r_u = %d",l_r_u);
	  #5 mem_resp = 1;
	  $display("initial l_r_u = %d",l_r_u);
	  #5 mem_resp = 0;
	  hit = 4'h4;
	  $display("initial l_r_u = %d",l_r_u);
	  #5 mem_resp = 1;
	  $display("initial l_r_u = %d",l_r_u);
	  #5 mem_resp = 0;
	  hit = 4'h8;
	  $display("initial l_r_u = %d",l_r_u);
	  #5 mem_resp = 1;
	  $display("initial l_r_u = %d",l_r_u);
	  #5 mem_resp = 0;
	  hit = 4'h1;
	  $display("initial l_r_u = %d",l_r_u);
	  #5 mem_resp = 1;
	  $display("initial l_r_u = %d",l_r_u);
	  #5 mem_resp = 0;
	  hit = 4'h2;
	  $display("initial l_r_u = %d",l_r_u);
	  #5 mem_resp = 1;
	  $display("initial l_r_u = %d",l_r_u);
	  #5 mem_resp = 0;
	  hit = 4'h4;
	  $display("initial l_r_u = %d",l_r_u);
	  #5 mem_resp = 1;
	  $display("initial l_r_u = %d",l_r_u);
	  #5 mem_resp = 0;
	  hit = 4'h8;
	  $display("initial l_r_u = %d",l_r_u);
	  #5 mem_resp = 1;
	  $display("initial l_r_u = %d",l_r_u);
	  #5 mem_resp = 0;
	  hit = 4'h0;
	  $display("initial l_r_u = %d",l_r_u);
	  #5 mem_resp = 1;
	  $display("initial l_r_u = %d",l_r_u);
	  #5 mem_resp = 0;
	  hit = 4'h4;
	  $display("initial l_r_u = %d",l_r_u);
	  #5 mem_resp = 1;
	  $display("initial l_r_u = %d",l_r_u);
	  #5 mem_resp = 0;
	  hit = 4'h2;
	  $display("initial l_r_u = %d",l_r_u);
	  #5 mem_resp = 1;
	  $display("initial l_r_u = %d",l_r_u);
	  #5 mem_resp = 0;
	  hit = 4'h2;
	  $display("initial l_r_u = %d",l_r_u);
	  #5 mem_resp = 1;
	  $display("initial l_r_u = %d",l_r_u);
	  #5 mem_resp = 0;
	  hit = 4'h1;
	  $display("l_r_u = %d",l_r_u);
	  #5 mem_resp=1;
	  $display("l_r_u = %d",l_r_u);

	  #5
	  hit = 4'h1;
	  mem_resp = 0;
	  $display("initial l_r_u = %d",l_r_u);
	  #5 mem_resp = 1;
	  $display("initial l_r_u = %d",l_r_u);
	  #5 mem_resp = 0;
	  hit = 4'h2;
	  $display("initial l_r_u = %d",l_r_u);
	  #5 mem_resp = 1;
	  $display("initial l_r_u = %d",l_r_u);
	  #5 mem_resp = 0;
	  hit = 4'h4;
	  $display("initial l_r_u = %d",l_r_u);
	  #5 mem_resp = 1;
	  $display("initial l_r_u = %d",l_r_u);
	  #5 mem_resp = 0;
	  hit = 4'h8;
	  $display("initial l_r_u = %d",l_r_u);
	  #5 mem_resp = 1;
	  $display("initial l_r_u = %d",l_r_u);
	  #5 mem_resp = 0;
	  hit = 4'h1;
	  $display("initial l_r_u = %d",l_r_u);
	  #5 mem_resp = 1;
	  $display("initial l_r_u = %d",l_r_u);
	  #5 mem_resp = 0;
	  hit = 4'h2;
	  $display("initial l_r_u = %d",l_r_u);
	  #5 mem_resp = 1;
	  $display("initial l_r_u = %d",l_r_u);
	  #5 mem_resp = 0;
	  hit = 4'h4;
	  $display("initial l_r_u = %d",l_r_u);
	  #5 mem_resp = 1;
	  $display("initial l_r_u = %d",l_r_u);
	  #5 mem_resp = 0;
	  hit = 4'h8;
	  $display("initial l_r_u = %d",l_r_u);
	  #5 mem_resp = 1;
	  $display("initial l_r_u = %d",l_r_u);
	  #5 mem_resp = 0;
	  hit = 4'h0;
	  $display("initial l_r_u = %d",l_r_u);
	  #5 mem_resp = 1;
	  $display("initial l_r_u = %d",l_r_u);
	  #5 mem_resp = 0;
	  hit = 4'h4;
	  $display("initial l_r_u = %d",l_r_u);
	  #5 mem_resp = 1;
	  $display("initial l_r_u = %d",l_r_u);
	  #5 mem_resp = 0;
	  hit = 4'h2;
	  $display("initial l_r_u = %d",l_r_u);
	  #5 mem_resp = 1;
	  $display("initial l_r_u = %d",l_r_u);
	  #5 mem_resp = 0;
	  hit = 4'h2;
	  $display("initial l_r_u = %d",l_r_u);
	  #5 mem_resp = 1;
	  $display("initial l_r_u = %d",l_r_u);
	  #5 mem_resp = 0;
	  hit = 4'h1;
	  $display("l_r_u = %d",l_r_u);
	  #5 mem_resp=1;
	  $display("l_r_u = %d",l_r_u);

	  #5
	  hit = 4'h1;
	  mem_resp = 0;
	  $display("initial l_r_u = %d",l_r_u);
	  #5 mem_resp = 1;
	  $display("initial l_r_u = %d",l_r_u);
	  #5 mem_resp = 0;
	  hit = 4'h2;
	  $display("initial l_r_u = %d",l_r_u);
	  #5 mem_resp = 1;
	  $display("initial l_r_u = %d",l_r_u);
	  #5 mem_resp = 0;
	  hit = 4'h4;
	  $display("initial l_r_u = %d",l_r_u);
	  #5 mem_resp = 1;
	  $display("initial l_r_u = %d",l_r_u);
	  #5 mem_resp = 0;
	  hit = 4'h8;
	  $display("initial l_r_u = %d",l_r_u);
	  #5 mem_resp = 1;
	  $display("initial l_r_u = %d",l_r_u);
	  #5 mem_resp = 0;
	  hit = 4'h1;
	  $display("initial l_r_u = %d",l_r_u);
	  #5 mem_resp = 1;
	  $display("initial l_r_u = %d",l_r_u);
	  #5 mem_resp = 0;
	  hit = 4'h2;
	  $display("initial l_r_u = %d",l_r_u);
	  #5 mem_resp = 1;
	  $display("initial l_r_u = %d",l_r_u);
	  #5 mem_resp = 0;
	  hit = 4'h4;
	  $display("initial l_r_u = %d",l_r_u);
	  #5 mem_resp = 1;
	  $display("initial l_r_u = %d",l_r_u);
	  #5 mem_resp = 0;
	  hit = 4'h8;
	  $display("initial l_r_u = %d",l_r_u);
	  #5 mem_resp = 1;
	  $display("initial l_r_u = %d",l_r_u);
	  #5 mem_resp = 0;
	  hit = 4'h0;
	  $display("initial l_r_u = %d",l_r_u);
	  #5 mem_resp = 1;
	  $display("initial l_r_u = %d",l_r_u);
	  #5 mem_resp = 0;
	  hit = 4'h4;
	  $display("initial l_r_u = %d",l_r_u);
	  #5 mem_resp = 1;
	  $display("initial l_r_u = %d",l_r_u);
	  #5 mem_resp = 0;
	  hit = 4'h2;
	  $display("initial l_r_u = %d",l_r_u);
	  #5 mem_resp = 1;
	  $display("initial l_r_u = %d",l_r_u);
	  #5 mem_resp = 0;
	  hit = 4'h2;
	  $display("initial l_r_u = %d",l_r_u);
	  #5 mem_resp = 1;
	  $display("initial l_r_u = %d",l_r_u);
	  #5 mem_resp = 0;
	  hit = 4'h1;
	  $display("l_r_u = %d",l_r_u);
	  #5 mem_resp=1;
	  $display("l_r_u = %d",l_r_u);

	  #5
	  hit = 4'h1;
	  mem_resp = 0;
	  $display("initial l_r_u = %d",l_r_u);
	  #5 mem_resp = 1;
	  $display("initial l_r_u = %d",l_r_u);
	  #5 mem_resp = 0;
	  hit = 4'h2;
	  $display("initial l_r_u = %d",l_r_u);
	  #5 mem_resp = 1;
	  $display("initial l_r_u = %d",l_r_u);
	  #5 mem_resp = 0;
	  hit = 4'h4;
	  $display("initial l_r_u = %d",l_r_u);
	  #5 mem_resp = 1;
	  $display("initial l_r_u = %d",l_r_u);
	  #5 mem_resp = 0;
	  hit = 4'h8;
	  $display("initial l_r_u = %d",l_r_u);
	  #5 mem_resp = 1;
	  $display("initial l_r_u = %d",l_r_u);
	  #5 mem_resp = 0;
	  hit = 4'h1;
	  $display("initial l_r_u = %d",l_r_u);
	  #5 mem_resp = 1;
	  $display("initial l_r_u = %d",l_r_u);
	  #5 mem_resp = 0;
	  hit = 4'h2;
	  $display("initial l_r_u = %d",l_r_u);
	  #5 mem_resp = 1;
	  $display("initial l_r_u = %d",l_r_u);
	  #5 mem_resp = 0;
	  hit = 4'h4;
	  $display("initial l_r_u = %d",l_r_u);
	  #5 mem_resp = 1;
	  $display("initial l_r_u = %d",l_r_u);
	  #5 mem_resp = 0;
	  hit = 4'h8;
	  $display("initial l_r_u = %d",l_r_u);
	  #5 mem_resp = 1;
	  $display("initial l_r_u = %d",l_r_u);
	  #5 mem_resp = 0;
	  hit = 4'h0;
	  $display("initial l_r_u = %d",l_r_u);
	  #5 mem_resp = 1;
	  $display("initial l_r_u = %d",l_r_u);
	  #5 mem_resp = 0;
	  hit = 4'h4;
	  $display("initial l_r_u = %d",l_r_u);
	  #5 mem_resp = 1;
	  $display("initial l_r_u = %d",l_r_u);
	  #5 mem_resp = 0;
	  hit = 4'h2;
	  $display("initial l_r_u = %d",l_r_u);
	  #5 mem_resp = 1;
	  $display("initial l_r_u = %d",l_r_u);
	  #5 mem_resp = 0;
	  hit = 4'h2;
	  $display("initial l_r_u = %d",l_r_u);
	  #5 mem_resp = 1;
	  $display("initial l_r_u = %d",l_r_u);
	  #5 mem_resp = 0;
	  hit = 4'h1;
	  $display("l_r_u = %d",l_r_u);
	  #5 mem_resp=1;
	  $display("l_r_u = %d",l_r_u);

	  #5
	  hit = 4'h1;
	  mem_resp = 0;
	  $display("initial l_r_u = %d",l_r_u);
	  #5 mem_resp = 1;
	  $display("initial l_r_u = %d",l_r_u);
	  #5 mem_resp = 0;
	  hit = 4'h2;
	  $display("initial l_r_u = %d",l_r_u);
	  #5 mem_resp = 1;
	  $display("initial l_r_u = %d",l_r_u);
	  #5 mem_resp = 0;
	  hit = 4'h4;
	  $display("initial l_r_u = %d",l_r_u);
	  #5 mem_resp = 1;
	  $display("initial l_r_u = %d",l_r_u);
	  #5 mem_resp = 0;
	  hit = 4'h8;
	  $display("initial l_r_u = %d",l_r_u);
	  #5 mem_resp = 1;
	  $display("initial l_r_u = %d",l_r_u);
	  #5 mem_resp = 0;
	  hit = 4'h1;
	  $display("initial l_r_u = %d",l_r_u);
	  #5 mem_resp = 1;
	  $display("initial l_r_u = %d",l_r_u);
	  #5 mem_resp = 0;
	  hit = 4'h2;
	  $display("initial l_r_u = %d",l_r_u);
	  #5 mem_resp = 1;
	  $display("initial l_r_u = %d",l_r_u);
	  #5 mem_resp = 0;
	  hit = 4'h4;
	  $display("initial l_r_u = %d",l_r_u);
	  #5 mem_resp = 1;
	  $display("initial l_r_u = %d",l_r_u);
	  #5 mem_resp = 0;
	  hit = 4'h8;
	  $display("initial l_r_u = %d",l_r_u);
	  #5 mem_resp = 1;
	  $display("initial l_r_u = %d",l_r_u);
	  #5 mem_resp = 0;
	  hit = 4'h0;
	  $display("initial l_r_u = %d",l_r_u);
	  #5 mem_resp = 1;
	  $display("initial l_r_u = %d",l_r_u);
	  #5 mem_resp = 0;
	  hit = 4'h4;
	  $display("initial l_r_u = %d",l_r_u);
	  #5 mem_resp = 1;
	  $display("initial l_r_u = %d",l_r_u);
	  #5 mem_resp = 0;
	  hit = 4'h2;
	  $display("initial l_r_u = %d",l_r_u);
	  #5 mem_resp = 1;
	  $display("initial l_r_u = %d",l_r_u);
	  #5 mem_resp = 0;
	  hit = 4'h2;
	  $display("initial l_r_u = %d",l_r_u);
	  #5 mem_resp = 1;
	  $display("initial l_r_u = %d",l_r_u);
	  #5 mem_resp = 0;
	  hit = 4'h1;
	  $display("l_r_u = %d",l_r_u);
	  #5 mem_resp=1;
	  $display("l_r_u = %d",l_r_u);

	  #5
	  hit = 4'h1;
	  mem_resp = 0;
	  $display("initial l_r_u = %d",l_r_u);
	  #5 mem_resp = 1;
	  $display("initial l_r_u = %d",l_r_u);
	  #5 mem_resp = 0;
	  hit = 4'h2;
	  $display("initial l_r_u = %d",l_r_u);
	  #5 mem_resp = 1;
	  $display("initial l_r_u = %d",l_r_u);
	  #5 mem_resp = 0;
	  hit = 4'h4;
	  $display("initial l_r_u = %d",l_r_u);
	  #5 mem_resp = 1;
	  $display("initial l_r_u = %d",l_r_u);
	  #5 mem_resp = 0;
	  hit = 4'h8;
	  $display("initial l_r_u = %d",l_r_u);
	  #5 mem_resp = 1;
	  $display("initial l_r_u = %d",l_r_u);
	  #5 mem_resp = 0;
	  hit = 4'h1;
	  $display("initial l_r_u = %d",l_r_u);
	  #5 mem_resp = 1;
	  $display("initial l_r_u = %d",l_r_u);
	  #5 mem_resp = 0;
	  hit = 4'h2;
	  $display("initial l_r_u = %d",l_r_u);
	  #5 mem_resp = 1;
	  $display("initial l_r_u = %d",l_r_u);
	  #5 mem_resp = 0;
	  hit = 4'h4;
	  $display("initial l_r_u = %d",l_r_u);
	  #5 mem_resp = 1;
	  $display("initial l_r_u = %d",l_r_u);
	  #5 mem_resp = 0;
	  hit = 4'h8;
	  $display("initial l_r_u = %d",l_r_u);
	  #5 mem_resp = 1;
	  $display("initial l_r_u = %d",l_r_u);
	  #5 mem_resp = 0;
	  hit = 4'h0;
	  $display("initial l_r_u = %d",l_r_u);
	  #5 mem_resp = 1;
	  $display("initial l_r_u = %d",l_r_u);
	  #5 mem_resp = 0;
	  hit = 4'h4;
	  $display("initial l_r_u = %d",l_r_u);
	  #5 mem_resp = 1;
	  $display("initial l_r_u = %d",l_r_u);
	  #5 mem_resp = 0;
	  hit = 4'h2;
	  $display("initial l_r_u = %d",l_r_u);
	  #5 mem_resp = 1;
	  $display("initial l_r_u = %d",l_r_u);
	  #5 mem_resp = 0;
	  hit = 4'h2;
	  $display("initial l_r_u = %d",l_r_u);
	  #5 mem_resp = 1;
	  $display("initial l_r_u = %d",l_r_u);
	  #5 mem_resp = 0;
	  hit = 4'h1;
	  $display("l_r_u = %d",l_r_u);
	  #5 mem_resp=1;
	  $display("l_r_u = %d",l_r_u);
   end : waveform_generation

endmodule // lru_tb
